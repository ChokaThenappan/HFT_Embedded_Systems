module avalon(
    input clk,
    input reset,
    input buffer_not_empty,
    input [7:0] ff_buffer_0,
    input [7:0] ff_buffer_1,
    input [7:0] ff_buffer_2,
    input [7:0] ff_buffer_3,
    input [7:0] ff_buffer_4,
    input [7:0] ff_buffer_5,
    input [7:0] ff_buffer_6,
    input [7:0] ff_buffer_7,
    input [7:0] ff_buffer_8,
    input [7:0] ff_buffer_9,
    input [7:0] ff_buffer_10,
    input [7:0] ff_buffer_11,
    input [7:0] ff_buffer_12,
    input [7:0] ff_buffer_13,
    input [7:0] ff_buffer_14,
    input [7:0] ff_buffer_15,
    input [7:0] ff_buffer_16,
    input [7:0] ff_buffer_17,
    input [7:0] ff_buffer_18,
    input [7:0] ff_buffer_19,
    input [7:0] ff_buffer_20,
    input [7:0] ff_buffer_21,
    input [7:0] ff_buffer_22,
    input [7:0] ff_buffer_23,
    input [7:0] ff_buffer_24,
    input [7:0] ff_buffer_25,
    input [7:0] ff_buffer_26,
    input [7:0] ff_buffer_27,
    input [7:0] ff_buffer_28,
    input [7:0] ff_buffer_29,
    input [7:0] ff_buffer_30,
    input [7:0] ff_buffer_31,
    input [7:0] ff_buffer_32,
    input [7:0] ff_buffer_33,
    input [7:0] ff_buffer_34,
    input [7:0] ff_buffer_35,
    input [7:0] ff_buffer_36,
    input [7:0] ff_buffer_37,
    input [7:0] ff_buffer_38,
    input [7:0] ff_buffer_39,
    input [7:0] ff_buffer_40,
    output logic system_free,
    output logic [7:0] max_order_id_1,
    output logic [7:0] max_quantity_1,
    output logic [7:0] max_price_1,
    output logic [7:0] max_order_id_2,
    output logic [7:0] max_quantity_2,
    output logic [7:0] max_price_2,
    output logic [7:0] max_order_id_3,
    output logic [7:0] max_quantity_3,
    output logic [7:0] max_price_3,
    output logic [7:0] max_order_id_4,
    output logic [7:0] max_quantity_4,
    output logic [7:0] max_price_4
);

top new_top (
    .clk(clk),
    .resetn(~reset),
    .buffer_not_empty(buffer_not_empty),
    .ff_buffer({ff_buffer_0, ff_buffer_1, ff_buffer_2, ff_buffer_3, ff_buffer_4, ff_buffer_5, ff_buffer_6, ff_buffer_7, ff_buffer_8, ff_buffer_9, ff_buffer_10, ff_buffer_11, ff_buffer_12, ff_buffer_13, ff_buffer_14, ff_buffer_15, ff_buffer_16, ff_buffer_17, ff_buffer_18, ff_buffer_19, ff_buffer_20, ff_buffer_21, ff_buffer_22, ff_buffer_23, ff_buffer_24, ff_buffer_25, ff_buffer_26, ff_buffer_27, ff_buffer_28, ff_buffer_29, ff_buffer_30, ff_buffer_31, ff_buffer_32, ff_buffer_33, ff_buffer_34, ff_buffer_35, ff_buffer_36, ff_buffer_37, ff_buffer_38, ff_buffer_39, ff_buffer_40}),
    .system_free(system_free),
    .max_order_id_1(max_order_id_1),
    .max_quantity_1(max_quantity_1),
    .max_price_1(max_price_1),
    .max_order_id_2(max_order_id_2),
    .max_quantity_2(max_quantity_2),
    .max_price_2(max_price_2),
    .max_order_id_3(max_order_id_3),
    .max_quantity_3(max_quantity_3),
    .max_price_3(max_price_3),
    .max_order_id_4(max_order_id_4),
    .max_quantity_4(max_quantity_4),
    .max_price_4(max_price_4)
);


endmodule
