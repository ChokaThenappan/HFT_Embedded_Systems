module avalon(
    input clk,
    input reset,
    input buffer_not_empty,
    input [31:0] ff_buffer_0,
    input [31:0] ff_buffer_1,
    input [31:0] ff_buffer_2,
    input [31:0] ff_buffer_3,
    input [31:0] ff_buffer_4,
    input [31:0] ff_buffer_5,
    input [31:0] ff_buffer_6,
    input [31:0] ff_buffer_7,
    input [31:0] ff_buffer_8,
    input [31:0] ff_buffer_9,
    input [31:0] ff_buffer_10,
    output logic system_free,
    output logic [31:0] max_order_id_1,
    output logic [31:0] max_quantity_1,
    output logic [31:0] max_price_1_1,
    output logic [31:0] max_price_1_2,
    output logic [31:0] max_order_id_2,
    output logic [31:0] max_quantity_2,
    output logic [31:0] max_price_2_1,
    output logic [31:0] max_price_2_2,
    output logic [31:0] max_order_id_3,
    output logic [31:0] max_quantity_3,
    output logic [31:0] max_price_3_1,
    output logic [31:0] max_price_3_2,
    output logic [31:0] max_order_id_4,
    output logic [31:0] max_quantity_4,
    output logic [31:0] max_price_4_1,
    output logic [31:0] max_price_4_2
);

top top_inst(
    .clk(clk),
    .resetn(~reset),
    .buffer_not_empty(buffer_not_empty),
    .ff_buffer({ff_buffer_0, ff_buffer_1, ff_buffer_2, ff_buffer_3, ff_buffer_4, ff_buffer_5, ff_buffer_6, ff_buffer_7, ff_buffer_8, ff_buffer_9, ff_buffer_10}),
    .system_free(system_free),
    .max_order_id_1(max_order_id_1),
    .max_quantity_1(max_quantity_1),
    .max_price_1({max_price_1_1, max_price_1_2}),
    .max_order_id_2(max_order_id_2),
    .max_quantity_2(max_quantity_2),
    .max_price_2({max_price_2_1, max_price_2_2}),
    .max_order_id_3(max_order_id_3),
    .max_quantity_3(max_quantity_3),
    .max_price_3({max_price_3_1, max_price_3_2}),
    .max_order_id_4(max_order_id_4),
    .max_quantity_4(max_quantity_4),
    .max_price_4({max_price_4_1, max_price_4_2})
);

endmodule
